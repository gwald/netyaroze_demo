pBAV       `� ��   @  ����Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������Sh@   ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    ��������  Sh    �������� @H        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   @N        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @N        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @\        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        ����� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����	 
 � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �  @dF       �����
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   8�||N..R\@	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      