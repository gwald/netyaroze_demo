pBAV        � ��   @  ����i�@   ��������i�@   ��������i�@   ��������i�@   ��������i�@   ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  i�    ��������  @H        �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ���\n�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    