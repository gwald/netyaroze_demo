pBAV       �[      @       �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             @@        ��               @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               Z=�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          