pBAV       � ��   @  ����d�	@   ���������	@   ���������	@   ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  �	    ��������  @H        �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   @7        �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @<      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   2.*�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        