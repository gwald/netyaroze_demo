pBAV       � ��q � N @  ����Z @   ��������Z @   ��������Z @   ��������Z @   ��������F @   ��������F @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������P @   ��������P @   ��������P @   ��������P @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������d @   ��������Z @   ��������Z @   ��������P @   ��������P @   ��������Z @   ��������n @   ��������n @   ��������n @   ��������n @   ��������d @   ��������d @   ��������d @   ��������d @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������d @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������_ @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������P @   ��������P @   ��������P @   ��������P @   ��������P @   ��������P @   ��������P @   ��������P @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������Z @   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       �������� @   �������� n@>& 5      ������   � � � �  @J 6A      ������   � � � �  @V'B      ����+�   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               �����_    � � � �               �����_    � � � �  n@>& A      ������  � � � �  @J BM      ������  � � � �  @V'N      ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  n@>& F      ������  � � � �  @J GR      ������  � � � �  @V'S      ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  Z@>& 5      ������  � � � �  k@J 6A      ������  � � � �  k@V'B      ����+�  � � � �  Z@> 5      ������  � � � �  k@J6A      ������  � � � �  k@VB      ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  @D| A      ����'�  � � � �  @P|B      ����'�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @D| A      ����'�  � � � �  @P|B      ����'�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @P| f      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  @P| f      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  @S: j    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @N> g      ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �  @S: j    ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �  @NF e    ����+� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @P|     ����+� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @P|     ����*�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @N> g      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @I| `    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Lm c    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Wy     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Wy     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Lm c    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @W~     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @W~     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @W~     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @W~     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @N* K    ������  � � � �  @N*Lc    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �  @N
 N    ������  � � � �  @N
Oe    ����'�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �  @B :    ����'�  � � � �  @N
;R    ������  � � � �  @N
Se    ����'�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @B ?    ����#�  � � � �  @N,@F    ������  � � � �  @N,Ge    ����#�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @K> b    ����%�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @1z 1    ������  � � � �  @={2=    ������  � � � �  @Iz>`    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  @1z 1    ������  � � � �  @={2=    ������  � � � �  @Iz>`    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �  @P{ g    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @/* E    ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   @#{ 9    ������!  � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �               ��    !   � � � �   @#{ 9    ������"  � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �               ��    "   � � � �   @#{ 9    ������#  � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �               ��    #   � � � �   @/, E    ������$  � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �               ��    $   � � � �   @/, E    ������%  � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �               ��    %   � � � �   @# 9    ������&  � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �               ��    &   � � � �   @# 9    ������'  � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �               ��    '   � � � �  @P| e    �����_(  � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �               ��    (   � � � �  @D| Z    �����)   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               ��    )   � � � �               �����_)   � � � �  @8| O    ������* ! � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               ��    *   � � � �               �����_*   � � � �  @8| O    ������+ ! � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               ��    +   � � � �               �����_+   � � � �  @T     ������, % � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               ��    ,   � � � �               �����_,   � � � �  @P$ d    ����,�- " � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �               ��    -   � � � �  @D| [    ������. # � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               ��    .   � � � �               �����_.   � � � �  @;n 4    ������/ $ � � � �  @;n5<    ����,�/ $ � � � �  @;n=J    ����+�/ $ � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �               ��    /   � � � �  @T     ������0 % � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               ��    0   � � � �               �����_0   � � � �  @T     ������1 % � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               ��    1   � � � �               �����_1   � � � �  @P e    ������2 & � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �               ��    2   � � � �  @P e    ������3 & � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �               ��    3   � � � �  @BB X    ��ק��4 ' � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               ��    4   � � � �               �����_4   � � � �  @BB X    ��ק��5 ' � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               ��    5   � � � �               �����_5   � � � �  n@BL X    ��ק��6 ' � � � �  n@B8 X    ��ק��6 ' � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               ��    6   � � � �               �����_6   � � � �  @XB i    ������7 ( � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �               ��    7   � � � �  @D| Y    ������8 ) � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �               �����_8   � � � �  @D| Y    ��؛��9 * � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �               �����_9   � � � �  @,| A    ��ڛ��: + � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �               �����_:   � � � �  @D| T    ������; , � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �               �����_;   � � � �  @G; [    ������< - � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �               �����_<   � � � �  @O8 d    ������= . � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �               �����_=   � � � �  @O# e    ������> / � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �               �����_>   � � � �  @O# e    ������? / � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �               �����_?   � � � �  @I| `    ������@ 0 � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �               �����_@   � � � �  @=| T    �����A 1 � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �               �����_A   � � � �  @=| T    ������B 2 � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �               �����_B   � � � �  @6| L    ������C 3 � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �               �����_C   � � � �  @P| e    ������D 4 � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �               �����_D   � � � �  @P|     ������E 5 � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �               �����_E   � � � �  @,| ,    ������F 6 � � � �  @8|-M    ������F 7 � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �               �����_F   � � � �  @I| `    ������G 8 � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �               �����_G   � � � �  @P| b    ������H 9 � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �               �����_H   � � � �  @P| R    ��ʩ��I : � � � �  @\|S    ��ʧ��I ; � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �               �����_I   � � � �  @P| e    ������J < � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �               �����_J   � � � �  @P| R    ��ʩ��K : � � � �  @\|S    ��ʧ��K ; � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �               �����_K   � � � �  @P| R    ��ʩ��L : � � � �  @\|S    ��ʧ��L ; � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �               �����_L   � � � �  w@NG e    ������M = � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �               �����_M   � � � �  @P| e    ������N < � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �               �����_N   � � � �  @P| e    ������O < � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �               �����_O   � � � �  @O# e    ������P / � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �               �����_P   � � � �  @O# e    ������Q / � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �               �����_Q   � � � �  @P| R    ��ʩ��R : � � � �  @\|S    ��ʧ��R ; � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �               �����_R   � � � �  @P| R    ��ʩ��S : � � � �  @\|S    ��ʧ��S ; � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �               �����_S   � � � �  @O# e    ������T / � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �               �����_T   � � � �  n@BL X    ��ק��U ' � � � �  n@B8 X    ��ק��U ' � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               ��    U   � � � �               �����_U   � � � �  @O# e    ������V / � � � �  n@T# e    ������V / � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �               �����_V   � � � �  @O# e    ������W / � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �               �����_W   � � � �  @ND d    �����X > � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �               �����_X   � � � �  @ND d    �����Y > � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �               �����_Y   � � � �  @ND d    �����Z > � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �               �����_Z   � � � �  @ND d    �����[ > � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �               �����_[   � � � �  @ND d    �����\ > � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �               �����_\   � � � �  @ND d    �����] > � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �               �����_]   � � � �  @ND d    �����^ > � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �               �����_^   � � � �  @ND d    �����_ > � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �               �����__   � � � �  @ND d    �����` > � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �               �����_`   � � � �  @ND d    �����a > � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �               �����_a   � � � �  @ND d    �����b > � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �               �����_b   � � � �  @ND d    �����c > � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �               �����_c   � � � �  @ND d    �����d > � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �               �����_d   � � � �  @ND d    �����e > � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �               �����_e   � � � �  @ND d    �����f > � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �               �����_f   � � � �  @ND d    �����g > � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �               �����_g   � � � �  @SG `    ����,�h ? � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �               �����_h   � � � �  @=| T    ������i @ � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �               �����_i   � � � �  @=| T    ������j @ � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �               �����_j   � � � �  @=| T    ����-�k A � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �               �����_k   � � � �  @P| e    ��d�-�l B � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �               �����_l   � � � �  @6| ;    ������m C � � � �  @P|<    ������m D � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �               �����_m   � � � �  @8| O    ������n ! � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               ��    n   � � � �               �����_n   � � � �  @D| Y    ������o E � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �               �����_o   � � � �   @-C#$      ������ F � � � �  n@+m%%      ������ G � � � �  @*F&&      ������ H � � � �  @+F''      ������ I � � � �  @*F((      ������ H � � � �  @C))      ������ K � � � �  @0F**      ����)� J � � � �  (=C++      ������ K � � � �  @2F,,      ����)� J � � � �  2;C--      ������ K � � � �  d@4F..      ������ J � � � �  @6C/0      ������ K � � � �  @?A11      ������ M � � � �  P2C22      ������ K � � � �  @9A33      ������ N � � � �  @>C55      ������ L � � � �   �z0�� >��f 6~ @(*J���$D`r (�`V� ,�T��t�l� �0\R�� (0� J � v � � � h � � 
R�*DL@ �� � ������n                                                                                                                                                                                                                                                                                                                                                                  